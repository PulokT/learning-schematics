* C:\Users\User\Desktop\New folder (2)\PSpice Solution for assignment 2  RL circuits only\RLRC updated\3RL.sch

* Schematics Version 9.2
* Wed Oct 23 02:37:52 2019



** Analysis setup **
.tran 0ns 122us 0ms 1us
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "3RL.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
